library verilog;
use verilog.vl_types.all;
entity compuerta_xor2_vlg_check_tst is
    port(
        SC              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end compuerta_xor2_vlg_check_tst;
