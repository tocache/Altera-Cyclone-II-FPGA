library verilog;
use verilog.vl_types.all;
entity xor_vhdl_vlg_check_tst is
    port(
        OUT_C           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end xor_vhdl_vlg_check_tst;
