library verilog;
use verilog.vl_types.all;
entity xor_vhdl_vlg_vec_tst is
end xor_vhdl_vlg_vec_tst;
