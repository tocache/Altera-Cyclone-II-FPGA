library verilog;
use verilog.vl_types.all;
entity el_ultimo_vlg_vec_tst is
end el_ultimo_vlg_vec_tst;
