library verilog;
use verilog.vl_types.all;
entity CKTO_4_vlg_check_tst is
    port(
        OD              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end CKTO_4_vlg_check_tst;
