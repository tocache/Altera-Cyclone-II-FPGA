library verilog;
use verilog.vl_types.all;
entity Compuerta_NAND_vlg_check_tst is
    port(
        OUTC            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Compuerta_NAND_vlg_check_tst;
