library verilog;
use verilog.vl_types.all;
entity CKTO_4_vlg_vec_tst is
end CKTO_4_vlg_vec_tst;
