library verilog;
use verilog.vl_types.all;
entity compuerta_xor_vlg_vec_tst is
end compuerta_xor_vlg_vec_tst;
