library verilog;
use verilog.vl_types.all;
entity nand_vhdl_vlg_vec_tst is
end nand_vhdl_vlg_vec_tst;
