library verilog;
use verilog.vl_types.all;
entity Compuerta_NAND_vlg_vec_tst is
end Compuerta_NAND_vlg_vec_tst;
