library verilog;
use verilog.vl_types.all;
entity ejemplo20211_1 is
    port(
        OUT_C           : out    vl_logic;
        IN_A            : in     vl_logic;
        IN_B            : in     vl_logic
    );
end ejemplo20211_1;
