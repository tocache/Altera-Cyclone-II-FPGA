library verilog;
use verilog.vl_types.all;
entity detect_vlg_vec_tst is
end detect_vlg_vec_tst;
