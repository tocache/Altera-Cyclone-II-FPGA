library verilog;
use verilog.vl_types.all;
entity Compuerta_XOR_vlg_vec_tst is
end Compuerta_XOR_vlg_vec_tst;
