library verilog;
use verilog.vl_types.all;
entity CKTO_3_vlg_vec_tst is
end CKTO_3_vlg_vec_tst;
