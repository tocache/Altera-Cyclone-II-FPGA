library verilog;
use verilog.vl_types.all;
entity \20211_el42_or1\ is
    port(
        OUT_C           : out    vl_logic;
        IN_B            : in     vl_logic;
        IN_A            : in     vl_logic
    );
end \20211_el42_or1\;
