library verilog;
use verilog.vl_types.all;
entity ejemplo20211_1_vlg_vec_tst is
end ejemplo20211_1_vlg_vec_tst;
