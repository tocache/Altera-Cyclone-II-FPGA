library verilog;
use verilog.vl_types.all;
entity compuerta_xor2_vlg_vec_tst is
end compuerta_xor2_vlg_vec_tst;
