library verilog;
use verilog.vl_types.all;
entity ejemplo20211_1_vlg_check_tst is
    port(
        OUT_C           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ejemplo20211_1_vlg_check_tst;
