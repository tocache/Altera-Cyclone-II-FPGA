library verilog;
use verilog.vl_types.all;
entity CKTO_3_vlg_check_tst is
    port(
        OUTD            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end CKTO_3_vlg_check_tst;
