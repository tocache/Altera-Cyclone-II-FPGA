library verilog;
use verilog.vl_types.all;
entity compuerta_xor_vlg_check_tst is
    port(
        OUT_C           : in     vl_logic;
        OUT_D           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end compuerta_xor_vlg_check_tst;
